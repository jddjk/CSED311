module immgen();

endmodule 
