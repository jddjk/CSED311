module alu_control_unit();

endmodule
