module add_alu (


);


endmodule