module pc();

endmodule
