module pc(
    input reset,
    input clk,
    input [31:0]next_pc,
    output reg [31:0]current_pc;
);

endmodule
